module wb_intercon
  #(parameter aw = 32,
    parameter dw = 32)
  (input 	   wb_clk_i,
   input 	   wb_rst_i,
   // OR1200 Instruction bus (To Master)
   input [aw-1:0]  wb_or1200_i_adr_i,
   input [dw-1:0]  wb_or1200_i_dat_i,
   input [3:0] 	   wb_or1200_i_sel_i,
   input 	   wb_or1200_i_we_i,
   input 	   wb_or1200_i_cyc_i,
   input 	   wb_or1200_i_stb_i,
   input [2:0] 	   wb_or1200_i_cti_i,
   input [1:0] 	   wb_or1200_i_bte_i,
   output [dw-1:0] wb_or1200_i_dat_o,
   output 	   wb_or1200_i_ack_o,
   output 	   wb_or1200_i_err_o,
   output 	   wb_or1200_i_rty_o,
   // OR1200 Data bus (To Master)
   input [aw-1:0]  wb_or1200_d_adr_i,
   input [dw-1:0]  wb_or1200_d_dat_i,
   input [3:0] 	   wb_or1200_d_sel_i,
   input 	   wb_or1200_d_we_i,
   input 	   wb_or1200_d_cyc_i,
   input 	   wb_or1200_d_stb_i,
   input [2:0] 	   wb_or1200_d_cti_i,
   input [1:0] 	   wb_or1200_d_bte_i,
   output [dw-1:0] wb_or1200_d_dat_o,
   output 	   wb_or1200_d_ack_o,
   output 	   wb_or1200_d_err_o,
   output 	   wb_or1200_d_rty_o,
   // Memory Interface (To Slave)
   output [aw-1:0] wb_mem_adr_o,
   output [dw-1:0] wb_mem_dat_o,
   output [3:0]    wb_mem_sel_o,
   output 	   wb_mem_we_o,
   output 	   wb_mem_cyc_o,
   output 	   wb_mem_stb_o,
   output [2:0]    wb_mem_cti_o,
   output [1:0]    wb_mem_bte_o,
   input [dw-1:0]  wb_mem_dat_i,
   input 	   wb_mem_ack_i,
   input 	   wb_mem_err_i,
   input 	   wb_mem_rty_i);

   //Memory Arbiter
   wb_arbiter wb_arbiter0
     (
      // Clock, reset
      .wb_clk_i				(wb_clk_i),
      .wb_rst_i				(wb_rst_i),
      // Wishbone slave interface 0
      .wbm0_adr_i			(wb_or1200_i_adr_i),
      .wbm0_dat_i			(wb_or1200_i_dat_i),
      .wbm0_sel_i			(wb_or1200_i_sel_i),
      .wbm0_we_i			(wb_or1200_i_we_i ),
      .wbm0_cyc_i			(wb_or1200_i_cyc_i),
      .wbm0_stb_i			(wb_or1200_i_stb_i),
      .wbm0_cti_i			(wb_or1200_i_cti_i),
      .wbm0_bte_i			(wb_or1200_i_bte_i),
      .wbm0_dat_o			(wb_or1200_i_dat_o),
      .wbm0_ack_o			(wb_or1200_i_ack_o),
      .wbm0_err_o                       (wb_or1200_i_err_o),
      .wbm0_rty_o                       (wb_or1200_i_rty_o),
      // Wishbone slave interface 1
      .wbm1_adr_i			(wb_or1200_d_adr_i),
      .wbm1_dat_i			(wb_or1200_d_dat_i),
      .wbm1_sel_i			(wb_or1200_d_sel_i),
      .wbm1_we_i			(wb_or1200_d_we_i),
      .wbm1_cyc_i			(wb_or1200_d_cyc_i),
      .wbm1_stb_i			(wb_or1200_d_stb_i),
      .wbm1_cti_i			(wb_or1200_d_cti_i),
      .wbm1_bte_i			(wb_or1200_d_bte_i),
      .wbm1_dat_o			(wb_or1200_d_dat_o),
      .wbm1_ack_o			(wb_or1200_d_ack_o),
      .wbm1_err_o                       (wb_or1200_d_err_o),
      .wbm1_rty_o                       (wb_or1200_d_rty_o),
      // Wishbone slave interface 2
      .wbm2_adr_i			(32'd0),
      .wbm2_dat_i			(32'd0),
      .wbm2_sel_i			(4'd0),
      .wbm2_cti_i			(3'd0),
      .wbm2_bte_i			(2'd0),
      .wbm2_we_i			(1'd0),
      .wbm2_cyc_i			(1'd0),
      .wbm2_stb_i			(1'd0),
      .wbm2_dat_o			(),
      .wbm2_ack_o			(),
      .wbm2_err_o                       (),
      .wbm2_rty_o                       (),
      //Wishbone Master interface
      .wbs_adr_o			(wb_mem_adr_o),
      .wbs_dat_o			(wb_mem_dat_o),
      .wbs_sel_o			(wb_mem_sel_o),
      .wbs_we_o			        (wb_mem_we_o ),
      .wbs_cyc_o			(wb_mem_cyc_o),
      .wbs_stb_o			(wb_mem_stb_o),
      .wbs_cti_o			(wb_mem_cti_o),
      .wbs_bte_o			(wb_mem_bte_o),
      .wbs_sdt_i			(wb_mem_dat_i),
      .wbs_ack_i			(wb_mem_ack_i),
      .wbs_err_i                        (wb_mem_err_i),
      .wbs_rty_i                        (wb_mem_rty_i));
         
endmodule // wb_intercon
